module Hazard2_SoC_tb;
    reg         HCLK;
    reg         HRESETn;

    wire [2:0] LED_out;

    
    // clock
    initial HCLK = 0;
    always #5 HCLK = ~HCLK;

    // Reset
    // initial begin
    //     HRESETn = 0;
    //     #47;
    //     @(posedge HCLK);
    //     HRESETn = 1;
    // end

    // TB infrastructure
    initial begin
        $dumpfile("Hazard2_SoC_tb.vcd");
        $dumpvars(0, Hazard2_SoC_tb);
        #10000;
        $display("Test Failed: Timeout");
        $finish;
    end

    Hazard2_SoC MUV (
        .HCLK(HCLK),
        // .HRESETn(HRESETn),
        .LED_out(LED_out)
    );




endmodule